<dec f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.h' l='65' type='QStringView'/>
<offset>256</offset>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='114' u='w' c='_ZN19QTextBoundaryFinderC1ERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='114' u='r' c='_ZN19QTextBoundaryFinderC1ERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='119' u='m' c='_ZN19QTextBoundaryFinderC1ERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='120' u='m' c='_ZN19QTextBoundaryFinderC1ERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='122' u='m' c='_ZN19QTextBoundaryFinderC1ERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='135' u='m' c='_ZN19QTextBoundaryFinderaSERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='136' u='m' c='_ZN19QTextBoundaryFinderaSERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='145' u='w' c='_ZN19QTextBoundaryFinderaSERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='145' u='r' c='_ZN19QTextBoundaryFinderaSERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='149' u='m' c='_ZN19QTextBoundaryFinderaSERKS_'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='175' u='w' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeERK7QString'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='180' u='m' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeERK7QString'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='181' u='m' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeERK7QString'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='183' u='r' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeERK7QString'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='210' u='w' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeE11QStringViewPhx'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='215' u='m' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeE11QStringViewPhx'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='216' u='m' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeE11QStringViewPhx'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='220' u='m' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeE11QStringViewPhx'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='223' u='r' c='_ZN19QTextBoundaryFinderC1ENS_12BoundaryTypeE11QStringViewPhx'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='244' u='m' c='_ZN19QTextBoundaryFinder5toEndEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='271' u='m' c='_ZN19QTextBoundaryFinder11setPositionEx'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='290' u='m' c='_ZNK19QTextBoundaryFinder6stringEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='290' u='m' c='_ZNK19QTextBoundaryFinder6stringEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='292' u='m' c='_ZNK19QTextBoundaryFinder6stringEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='303' u='m' c='_ZN19QTextBoundaryFinder14toNextBoundaryEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='311' u='m' c='_ZN19QTextBoundaryFinder14toNextBoundaryEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='315' u='m' c='_ZN19QTextBoundaryFinder14toNextBoundaryEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='319' u='m' c='_ZN19QTextBoundaryFinder14toNextBoundaryEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='323' u='m' c='_ZN19QTextBoundaryFinder14toNextBoundaryEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='338' u='m' c='_ZN19QTextBoundaryFinder18toPreviousBoundaryEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='371' u='m' c='_ZNK19QTextBoundaryFinder12isAtBoundaryEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='394' u='m' c='_ZNK19QTextBoundaryFinder15boundaryReasonsEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='404' u='m' c='_ZNK19QTextBoundaryFinder15boundaryReasonsEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='422' u='m' c='_ZNK19QTextBoundaryFinder15boundaryReasonsEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='434' u='m' c='_ZNK19QTextBoundaryFinder15boundaryReasonsEv'/>
<use f='qtbase-6.5.0/src/corelib/text/qtextboundaryfinder.cpp' l='436' u='m' c='_ZNK19QTextBoundaryFinder15boundaryReasonsEv'/>
