<dec f='qtbase-6.5.0/src/gui/painting/qpainter_p.h' l='133' type='int'/>
<offset>3232</offset>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='211' u='r' c='_ZNK15QPainterPrivate13viewTransformEv'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='264' u='w' c='_ZN15QPainterPrivate20attachPainterPrivateEP8QPainterP12QPaintDevice'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='1786' u='w' c='_ZN8QPainter5beginEP12QPaintDevice'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='1816' u='w' c='_ZN8QPainter5beginEP12QPaintDevice'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='1819' u='w' c='_ZN8QPainter5beginEP12QPaintDevice'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='7015' u='w' c='_ZN8QPainter11setViewportERK5QRect'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='7034' u='r' c='_ZNK8QPainter8viewportEv'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='7357' u='w' c='_ZN13QPainterStateC1EPKS_'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='7357' u='r' c='_ZN13QPainterStateC1EPKS_'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='7384' u='w' c='_ZN13QPainterState4initEP8QPainter'/>
<use f='qtbase-6.5.0/src/gui/painting/qpainter.cpp' l='7903' u='w' c='_ZN8QPainter14resetTransformEv'/>
